module ConstMemory( Data , Address , WriteEnable , Clock , Reset );
    parameter           Size    =   256;
    
    inout  [47:0]       Data;
    input  [ 7:0]       Address;
    input               WriteEnable;
    input               Clock;
    input               Reset;
    
    reg  [47:0]         Memory[Size-1:0];
    
    wire [47:0]         ip;
    wire [47:0]         op;
    
    bufif1              b1[47:0]    ( Data , op   , ~WriteEnable );
    bufif1              b2[47:0]    ( ip   , Data ,  WriteEnable );
    
    assign  op          =   Memory[Address];
    
    always @(negedge Reset , posedge Clock)
    begin
        if(!Reset)
        begin
            Memory[0]     <=  48'h8000_4000_0000;       //  2 v0 +          // 2 v0 + 11 v4 ;   44
            Memory[1]     <=  48'h8001_4040_0000;       //  3 v1 +          // 3 v1 + 13 v5;    -62
            Memory[2]     <=  48'hC002_40A0_0000;       //  5 v2 ;  10
            Memory[3]     <=  48'hC003_40E0_0000;       //  7 v3 ;  21
            Memory[4]     <=  48'h4004_4130_0000;       // + 11 v4 ;        //  2 v1 + 11 v4;
            Memory[5]     <=  48'h4005_4150_0000;       // + 13 v5 +        //  3 v2 + 13 v5 ;
            Memory[6]     <=  48'h0000_0000_0000;       
            Memory[7]     <=  48'h0000_0000_0000;       // xxx
            Memory[8]     <=  48'h0000_0000_0000;       // xxx
            Memory[9]     <=  48'h2000_0000_0000;       // + 17 v8 ;        //  3 v2 + 13 v6 + 17 v8 ;
            Memory[10]    <=  48'h0000_0000_0000;       // + 19 v9 ;        // 16 v7 + 19 v9 ;
            Memory[11]    <=  48'h0000_0000_0000;       // xxx
            Memory[12]    <=  48'h0000_0000_0000;
            Memory[13]    <=  48'h0000_0000_0000;
            Memory[14]    <=  48'h2000_0000_0000;       // End-of-all-equations bit
            Memory[15]    <=  48'h0000_0000_0000;
            Memory[16]    <=  48'h0000_0000_0000;       // + 11 v5 ;        //  2 v1 + 11 v5 ;
            Memory[17]    <=  48'h0000_0000_0000;       // + 13 v6 +        //  3 v2 + 13 v6 + 17 v8 ;
            Memory[18]    <=  48'h0000_0000_0000;       //   16 v7 +        // 16 v7 + 19 v9 ;
            Memory[19]    <=  48'h0000_0000_0000;       // xxx
            Memory[20]    <=  48'h0000_0000_0000;
            Memory[21]    <=  48'h0000_0000_0000;
            Memory[22]    <=  48'h0000_0000_0000;
            Memory[23]    <=  48'h0000_0000_0000;
            Memory[24]    <=  48'h0000_0000_0000;
            Memory[25]    <=  48'h0000_0000_0000;
            Memory[26]    <=  48'h0000_0000_0000;
            Memory[27]    <=  48'h0000_0000_0000;
            Memory[28]    <=  48'h0000_0000_0000;
            Memory[29]    <=  48'h0000_0000_0000;
            Memory[30]    <=  48'h0000_0000_0000;
            Memory[31]    <=  48'h0000_0000_0000;
            Memory[32]    <=  48'h0000_0000_0000;       // xxx
            Memory[33]    <=  48'h4008_4188_0000;       // + 17 v8 ;        //  3 v2 + 13 v6 + 17 v8 ;
            Memory[34]    <=  48'h4009_4198_0000;       // + 19 v9 ;        // 16 v7 + 19 v9 ;
            Memory[35]    <=  48'h0000_0000_0000;       // xxx
            Memory[36]    <=  48'h0000_0000_0000;
            Memory[37]    <=  48'h0000_0000_0000;
            Memory[38]    <=  48'h0000_0000_0000;
            Memory[39]    <=  48'h0000_0000_0000;
            Memory[40]    <=  48'h0000_0000_0000;
            Memory[41]    <=  48'h0000_0000_0000;
            Memory[42]    <=  48'h0000_0000_0000;
            Memory[43]    <=  48'h0000_0000_0000;
            Memory[44]    <=  48'h0000_0000_0000;
            Memory[45]    <=  48'h0000_0000_0000;
            Memory[46]    <=  48'h0000_0000_0000;
            Memory[47]    <=  48'h0000_0000_0000;
            Memory[48]    <=  48'h0000_0000_0000;
            Memory[49]    <=  48'h0000_0000_0000;
            Memory[50]    <=  48'h2000_0000_0000;       // Stall bit
            Memory[51]    <=  48'h0000_0000_0000;
            Memory[52]    <=  48'h0000_0000_0000;
            Memory[53]    <=  48'h0000_0000_0000;
            Memory[54]    <=  48'h0000_0000_0000;
            Memory[55]    <=  48'h0000_0000_0000;
            Memory[56]    <=  48'h0000_0000_0000;
            Memory[57]    <=  48'h0000_0000_0000;
            Memory[58]    <=  48'h0000_0000_0000;
            Memory[59]    <=  48'h0000_0000_0000;
            Memory[60]    <=  48'h0000_0000_0000;
            Memory[61]    <=  48'h0000_0000_0000;
            Memory[62]    <=  48'h0000_0000_0000;
            Memory[63]    <=  48'h0000_0000_0000;
            Memory[64]    <=  48'h0000_0000_0000;
            Memory[65]    <=  48'h0000_0000_0000;
            Memory[66]    <=  48'h0000_0000_0000;
            Memory[67]    <=  48'h0000_0000_0000;
            Memory[68]    <=  48'h0000_0000_0000;
            Memory[69]    <=  48'h0000_0000_0000;
            Memory[70]    <=  48'h0000_0000_0000;
            Memory[71]    <=  48'h0000_0000_0000;
            Memory[72]    <=  48'h0000_0000_0000;
            Memory[73]    <=  48'h0000_0000_0000;
            Memory[74]    <=  48'h0000_0000_0000;
            Memory[75]    <=  48'h0000_0000_0000;
            Memory[76]    <=  48'h0000_0000_0000;
            Memory[77]    <=  48'h0000_0000_0000;
            Memory[78]    <=  48'h0000_0000_0000;
            Memory[79]    <=  48'h0000_0000_0000;
            Memory[80]    <=  48'h0000_0000_0000;
            Memory[81]    <=  48'h0000_0000_0000;
            Memory[82]    <=  48'h0000_0000_0000;
            Memory[83]    <=  48'h0000_0000_0000;
            Memory[84]    <=  48'h0000_0000_0000;
            Memory[85]    <=  48'h0000_0000_0000;
            Memory[86]    <=  48'h0000_0000_0000;
            Memory[87]    <=  48'h0000_0000_0000;
            Memory[88]    <=  48'h0000_0000_0000;
            Memory[89]    <=  48'h0000_0000_0000;
            Memory[90]    <=  48'h0000_0000_0000;
            Memory[91]    <=  48'h0000_0000_0000;
            Memory[92]    <=  48'h0000_0000_0000;
            Memory[93]    <=  48'h0000_0000_0000;
            Memory[94]    <=  48'h0000_0000_0000;
            Memory[95]    <=  48'h0000_0000_0000;
            Memory[96]    <=  48'h0000_0000_0000;
            Memory[97]    <=  48'h0000_0000_0000;
            Memory[98]    <=  48'h0000_0000_0000;
            Memory[99]    <=  48'h0000_0000_0000;
            Memory[100]   <=  48'h0000_0000_0000;
            Memory[101]   <=  48'h0000_0000_0000;
            Memory[102]   <=  48'h0000_0000_0000;
            Memory[103]   <=  48'h0000_0000_0000;
            Memory[104]   <=  48'h0000_0000_0000;
            Memory[105]   <=  48'h0000_0000_0000;
            Memory[106]   <=  48'h0000_0000_0000;
            Memory[107]   <=  48'h0000_0000_0000;
            Memory[108]   <=  48'h0000_0000_0000;
            Memory[109]   <=  48'h0000_0000_0000;
            Memory[110]   <=  48'h0000_0000_0000;
            Memory[111]   <=  48'h0000_0000_0000;
            Memory[112]   <=  48'h0000_0000_0000;
            Memory[113]   <=  48'h0000_0000_0000;
            Memory[114]   <=  48'h0000_0000_0000;
            Memory[115]   <=  48'h0000_0000_0000;
            Memory[116]   <=  48'h0000_0000_0000;
            Memory[117]   <=  48'h0000_0000_0000;
            Memory[118]   <=  48'h0000_0000_0000;
            Memory[119]   <=  48'h0000_0000_0000;
            Memory[120]   <=  48'h0000_0000_0000;
            Memory[121]   <=  48'h0000_0000_0000;
            Memory[122]   <=  48'h0000_0000_0000;
            Memory[123]   <=  48'h0000_0000_0000;
            Memory[124]   <=  48'h0000_0000_0000;
            Memory[125]   <=  48'h0000_0000_0000;
            Memory[126]   <=  48'h0000_0000_0000;
            Memory[127]   <=  48'h0000_0000_0000;
            Memory[128]   <=  48'h0000_0000_0000;
            Memory[129]   <=  48'h0000_0000_0000;
            Memory[130]   <=  48'h0000_0000_0000;
            Memory[131]   <=  48'h0000_0000_0000;
            Memory[132]   <=  48'h0000_0000_0000;
            Memory[133]   <=  48'h0000_0000_0000;
            Memory[134]   <=  48'h0000_0000_0000;
            Memory[135]   <=  48'h0000_0000_0000;
            Memory[136]   <=  48'h0000_0000_0000;
            Memory[137]   <=  48'h0000_0000_0000;
            Memory[138]   <=  48'h0000_0000_0000;
            Memory[139]   <=  48'h0000_0000_0000;
            Memory[140]   <=  48'h0000_0000_0000;
            Memory[141]   <=  48'h0000_0000_0000;
            Memory[142]   <=  48'h0000_0000_0000;
            Memory[143]   <=  48'h0000_0000_0000;
            Memory[144]   <=  48'h0000_0000_0000;
            Memory[145]   <=  48'h0000_0000_0000;
            Memory[146]   <=  48'h0000_0000_0000;
            Memory[147]   <=  48'h0000_0000_0000;
            Memory[148]   <=  48'h0000_0000_0000;
            Memory[149]   <=  48'h0000_0000_0000;
            Memory[150]   <=  48'h0000_0000_0000;
            Memory[151]   <=  48'h0000_0000_0000;
            Memory[152]   <=  48'h0000_0000_0000;
            Memory[153]   <=  48'h0000_0000_0000;
            Memory[154]   <=  48'h0000_0000_0000;
            Memory[155]   <=  48'h0000_0000_0000;
            Memory[156]   <=  48'h0000_0000_0000;
            Memory[157]   <=  48'h0000_0000_0000;
            Memory[158]   <=  48'h0000_0000_0000;
            Memory[159]   <=  48'h0000_0000_0000;
            Memory[160]   <=  48'h0000_0000_0000;
            Memory[161]   <=  48'h0000_0000_0000;
            Memory[162]   <=  48'h0000_0000_0000;
            Memory[163]   <=  48'h0000_0000_0000;
            Memory[164]   <=  48'h0000_0000_0000;
            Memory[165]   <=  48'h0000_0000_0000;
            Memory[166]   <=  48'h0000_0000_0000;
            Memory[167]   <=  48'h0000_0000_0000;
            Memory[168]   <=  48'h0000_0000_0000;
            Memory[169]   <=  48'h0000_0000_0000;
            Memory[170]   <=  48'h0000_0000_0000;
            Memory[171]   <=  48'h0000_0000_0000;
            Memory[172]   <=  48'h0000_0000_0000;
            Memory[173]   <=  48'h0000_0000_0000;
            Memory[174]   <=  48'h0000_0000_0000;
            Memory[175]   <=  48'h0000_0000_0000;
            Memory[176]   <=  48'h0000_0000_0000;
            Memory[177]   <=  48'h0000_0000_0000;
            Memory[178]   <=  48'h0000_0000_0000;
            Memory[179]   <=  48'h0000_0000_0000;
            Memory[180]   <=  48'h0000_0000_0000;
            Memory[181]   <=  48'h0000_0000_0000;
            Memory[182]   <=  48'h0000_0000_0000;
            Memory[183]   <=  48'h0000_0000_0000;
            Memory[184]   <=  48'h0000_0000_0000;
            Memory[185]   <=  48'h0000_0000_0000;
            Memory[186]   <=  48'h0000_0000_0000;
            Memory[187]   <=  48'h0000_0000_0000;
            Memory[188]   <=  48'h0000_0000_0000;
            Memory[189]   <=  48'h0000_0000_0000;
            Memory[190]   <=  48'h0000_0000_0000;
            Memory[191]   <=  48'h0000_0000_0000;
            Memory[192]   <=  48'h0000_0000_0000;
            Memory[193]   <=  48'h0000_0000_0000;
            Memory[194]   <=  48'h0000_0000_0000;
            Memory[195]   <=  48'h0000_0000_0000;
            Memory[196]   <=  48'h0000_0000_0000;
            Memory[197]   <=  48'h0000_0000_0000;
            Memory[198]   <=  48'h0000_0000_0000;
            Memory[199]   <=  48'h0000_0000_0000;
            Memory[200]   <=  48'h0000_0000_0000;
            Memory[201]   <=  48'h0000_0000_0000;
            Memory[202]   <=  48'h0000_0000_0000;
            Memory[203]   <=  48'h0000_0000_0000;
            Memory[204]   <=  48'h0000_0000_0000;
            Memory[205]   <=  48'h0000_0000_0000;
            Memory[206]   <=  48'h0000_0000_0000;
            Memory[207]   <=  48'h0000_0000_0000;
            Memory[208]   <=  48'h0000_0000_0000;
            Memory[209]   <=  48'h0000_0000_0000;
            Memory[210]   <=  48'h0000_0000_0000;
            Memory[211]   <=  48'h0000_0000_0000;
            Memory[212]   <=  48'h0000_0000_0000;
            Memory[213]   <=  48'h0000_0000_0000;
            Memory[214]   <=  48'h0000_0000_0000;
            Memory[215]   <=  48'h0000_0000_0000;
            Memory[216]   <=  48'h0000_0000_0000;
            Memory[217]   <=  48'h0000_0000_0000;
            Memory[218]   <=  48'h0000_0000_0000;
            Memory[219]   <=  48'h0000_0000_0000;
            Memory[220]   <=  48'h0000_0000_0000;
            Memory[221]   <=  48'h0000_0000_0000;
            Memory[222]   <=  48'h0000_0000_0000;
            Memory[223]   <=  48'h0000_0000_0000;
            Memory[224]   <=  48'h0000_0000_0000;
            Memory[225]   <=  48'h0000_0000_0000;
            Memory[226]   <=  48'h0000_0000_0000;
            Memory[227]   <=  48'h0000_0000_0000;
            Memory[228]   <=  48'h0000_0000_0000;
            Memory[229]   <=  48'h0000_0000_0000;
            Memory[230]   <=  48'h0000_0000_0000;
            Memory[231]   <=  48'h0000_0000_0000;
            Memory[232]   <=  48'h0000_0000_0000;
            Memory[233]   <=  48'h0000_0000_0000;
            Memory[234]   <=  48'h0000_0000_0000;
            Memory[235]   <=  48'h0000_0000_0000;
            Memory[236]   <=  48'h0000_0000_0000;
            Memory[237]   <=  48'h0000_0000_0000;
            Memory[238]   <=  48'h0000_0000_0000;
            Memory[239]   <=  48'h0000_0000_0000;
            Memory[240]   <=  48'h0000_0000_0000;
            Memory[241]   <=  48'h0000_0000_0000;
            Memory[242]   <=  48'h0000_0000_0000;
            Memory[243]   <=  48'h0000_0000_0000;
            Memory[244]   <=  48'h0000_0000_0000;
            Memory[245]   <=  48'h0000_0000_0000;
            Memory[246]   <=  48'h0000_0000_0000;
            Memory[247]   <=  48'h0000_0000_0000;
            Memory[248]   <=  48'h0000_0000_0000;
            Memory[249]   <=  48'h0000_0000_0000;
            Memory[250]   <=  48'h0000_0000_0000;
            Memory[251]   <=  48'h0000_0000_0000;
            Memory[252]   <=  48'h0000_0000_0000;
            Memory[253]   <=  48'h0000_0000_0000;
            Memory[254]   <=  48'h0000_0000_0000;
            Memory[255]   <=  48'h0000_0000_0000;
        end
        else
        begin
            if(WriteEnable)
            begin
                Memory[Address] <=  ip;
            end
            else
            begin
                Memory[0]     <=  Memory[0];
                Memory[1]     <=  Memory[1];
                Memory[2]     <=  Memory[2];
                Memory[3]     <=  Memory[3];
                Memory[4]     <=  Memory[4];
                Memory[5]     <=  Memory[5];
                Memory[6]     <=  Memory[6];
                Memory[7]     <=  Memory[7];
                Memory[8]     <=  Memory[8];
                Memory[9]     <=  Memory[9];
                Memory[10]    <=  Memory[10];
                Memory[11]    <=  Memory[11];
                Memory[12]    <=  Memory[12];
                Memory[13]    <=  Memory[13];
                Memory[14]    <=  Memory[14];
                Memory[15]    <=  Memory[15];
                Memory[16]    <=  Memory[16];
                Memory[17]    <=  Memory[17];
                Memory[18]    <=  Memory[18];
                Memory[19]    <=  Memory[19];
                Memory[20]    <=  Memory[20];
                Memory[21]    <=  Memory[21];
                Memory[22]    <=  Memory[22];
                Memory[23]    <=  Memory[23];
                Memory[24]    <=  Memory[24];
                Memory[25]    <=  Memory[25];
                Memory[26]    <=  Memory[26];
                Memory[27]    <=  Memory[27];
                Memory[28]    <=  Memory[28];
                Memory[29]    <=  Memory[29];
                Memory[30]    <=  Memory[30];
                Memory[31]    <=  Memory[31];
                Memory[32]    <=  Memory[32];
                Memory[33]    <=  Memory[33];
                Memory[34]    <=  Memory[34];
                Memory[35]    <=  Memory[35];
                Memory[36]    <=  Memory[36];
                Memory[37]    <=  Memory[37];
                Memory[38]    <=  Memory[38];
                Memory[39]    <=  Memory[39];
                Memory[40]    <=  Memory[40];
                Memory[41]    <=  Memory[41];
                Memory[42]    <=  Memory[42];
                Memory[43]    <=  Memory[43];
                Memory[44]    <=  Memory[44];
                Memory[45]    <=  Memory[45];
                Memory[46]    <=  Memory[46];
                Memory[47]    <=  Memory[47];
                Memory[48]    <=  Memory[48];
                Memory[49]    <=  Memory[49];
                Memory[50]    <=  Memory[50];
                Memory[51]    <=  Memory[51];
                Memory[52]    <=  Memory[52];
                Memory[53]    <=  Memory[53];
                Memory[54]    <=  Memory[54];
                Memory[55]    <=  Memory[55];
                Memory[56]    <=  Memory[56];
                Memory[57]    <=  Memory[57];
                Memory[58]    <=  Memory[58];
                Memory[59]    <=  Memory[59];
                Memory[60]    <=  Memory[60];
                Memory[61]    <=  Memory[61];
                Memory[62]    <=  Memory[62];
                Memory[63]    <=  Memory[63];
                Memory[64]    <=  Memory[64];
                Memory[65]    <=  Memory[65];
                Memory[66]    <=  Memory[66];
                Memory[67]    <=  Memory[67];
                Memory[68]    <=  Memory[68];
                Memory[69]    <=  Memory[69];
                Memory[70]    <=  Memory[70];
                Memory[71]    <=  Memory[71];
                Memory[72]    <=  Memory[72];
                Memory[73]    <=  Memory[73];
                Memory[74]    <=  Memory[74];
                Memory[75]    <=  Memory[75];
                Memory[76]    <=  Memory[76];
                Memory[77]    <=  Memory[77];
                Memory[78]    <=  Memory[78];
                Memory[79]    <=  Memory[79];
                Memory[80]    <=  Memory[80];
                Memory[81]    <=  Memory[81];
                Memory[82]    <=  Memory[82];
                Memory[83]    <=  Memory[83];
                Memory[84]    <=  Memory[84];
                Memory[85]    <=  Memory[85];
                Memory[86]    <=  Memory[86];
                Memory[87]    <=  Memory[87];
                Memory[88]    <=  Memory[88];
                Memory[89]    <=  Memory[89];
                Memory[90]    <=  Memory[90];
                Memory[91]    <=  Memory[91];
                Memory[92]    <=  Memory[92];
                Memory[93]    <=  Memory[93];
                Memory[94]    <=  Memory[94];
                Memory[95]    <=  Memory[95];
                Memory[96]    <=  Memory[96];
                Memory[97]    <=  Memory[97];
                Memory[98]    <=  Memory[98];
                Memory[99]    <=  Memory[99];
                Memory[100]   <=  Memory[100];
                Memory[101]   <=  Memory[101];
                Memory[102]   <=  Memory[102];
                Memory[103]   <=  Memory[103];
                Memory[104]   <=  Memory[104];
                Memory[105]   <=  Memory[105];
                Memory[106]   <=  Memory[106];
                Memory[107]   <=  Memory[107];
                Memory[108]   <=  Memory[108];
                Memory[109]   <=  Memory[109];
                Memory[110]   <=  Memory[110];
                Memory[111]   <=  Memory[111];
                Memory[112]   <=  Memory[112];
                Memory[113]   <=  Memory[113];
                Memory[114]   <=  Memory[114];
                Memory[115]   <=  Memory[115];
                Memory[116]   <=  Memory[116];
                Memory[117]   <=  Memory[117];
                Memory[118]   <=  Memory[118];
                Memory[119]   <=  Memory[119];
                Memory[120]   <=  Memory[120];
                Memory[121]   <=  Memory[121];
                Memory[122]   <=  Memory[122];
                Memory[123]   <=  Memory[123];
                Memory[124]   <=  Memory[124];
                Memory[125]   <=  Memory[125];
                Memory[126]   <=  Memory[126];
                Memory[127]   <=  Memory[127];
                Memory[128]   <=  Memory[128];
                Memory[129]   <=  Memory[129];
                Memory[130]   <=  Memory[130];
                Memory[131]   <=  Memory[131];
                Memory[132]   <=  Memory[132];
                Memory[133]   <=  Memory[133];
                Memory[134]   <=  Memory[134];
                Memory[135]   <=  Memory[135];
                Memory[136]   <=  Memory[136];
                Memory[137]   <=  Memory[137];
                Memory[138]   <=  Memory[138];
                Memory[139]   <=  Memory[139];
                Memory[140]   <=  Memory[140];
                Memory[141]   <=  Memory[141];
                Memory[142]   <=  Memory[142];
                Memory[143]   <=  Memory[143];
                Memory[144]   <=  Memory[144];
                Memory[145]   <=  Memory[145];
                Memory[146]   <=  Memory[146];
                Memory[147]   <=  Memory[147];
                Memory[148]   <=  Memory[148];
                Memory[149]   <=  Memory[149];
                Memory[150]   <=  Memory[150];
                Memory[151]   <=  Memory[151];
                Memory[152]   <=  Memory[152];
                Memory[153]   <=  Memory[153];
                Memory[154]   <=  Memory[154];
                Memory[155]   <=  Memory[155];
                Memory[156]   <=  Memory[156];
                Memory[157]   <=  Memory[157];
                Memory[158]   <=  Memory[158];
                Memory[159]   <=  Memory[159];
                Memory[160]   <=  Memory[160];
                Memory[161]   <=  Memory[161];
                Memory[162]   <=  Memory[162];
                Memory[163]   <=  Memory[163];
                Memory[164]   <=  Memory[164];
                Memory[165]   <=  Memory[165];
                Memory[166]   <=  Memory[166];
                Memory[167]   <=  Memory[167];
                Memory[168]   <=  Memory[168];
                Memory[169]   <=  Memory[169];
                Memory[170]   <=  Memory[170];
                Memory[171]   <=  Memory[171];
                Memory[172]   <=  Memory[172];
                Memory[173]   <=  Memory[173];
                Memory[174]   <=  Memory[174];
                Memory[175]   <=  Memory[175];
                Memory[176]   <=  Memory[176];
                Memory[177]   <=  Memory[177];
                Memory[178]   <=  Memory[178];
                Memory[179]   <=  Memory[179];
                Memory[180]   <=  Memory[180];
                Memory[181]   <=  Memory[181];
                Memory[182]   <=  Memory[182];
                Memory[183]   <=  Memory[183];
                Memory[184]   <=  Memory[184];
                Memory[185]   <=  Memory[185];
                Memory[186]   <=  Memory[186];
                Memory[187]   <=  Memory[187];
                Memory[188]   <=  Memory[188];
                Memory[189]   <=  Memory[189];
                Memory[190]   <=  Memory[190];
                Memory[191]   <=  Memory[191];
                Memory[192]   <=  Memory[192];
                Memory[193]   <=  Memory[193];
                Memory[194]   <=  Memory[194];
                Memory[195]   <=  Memory[195];
                Memory[196]   <=  Memory[196];
                Memory[197]   <=  Memory[197];
                Memory[198]   <=  Memory[198];
                Memory[199]   <=  Memory[199];
                Memory[200]   <=  Memory[200];
                Memory[201]   <=  Memory[201];
                Memory[202]   <=  Memory[202];
                Memory[203]   <=  Memory[203];
                Memory[204]   <=  Memory[204];
                Memory[205]   <=  Memory[205];
                Memory[206]   <=  Memory[206];
                Memory[207]   <=  Memory[207];
                Memory[208]   <=  Memory[208];
                Memory[209]   <=  Memory[209];
                Memory[210]   <=  Memory[210];
                Memory[211]   <=  Memory[211];
                Memory[212]   <=  Memory[212];
                Memory[213]   <=  Memory[213];
                Memory[214]   <=  Memory[214];
                Memory[215]   <=  Memory[215];
                Memory[216]   <=  Memory[216];
                Memory[217]   <=  Memory[217];
                Memory[218]   <=  Memory[218];
                Memory[219]   <=  Memory[219];
                Memory[220]   <=  Memory[220];
                Memory[221]   <=  Memory[221];
                Memory[222]   <=  Memory[222];
                Memory[223]   <=  Memory[223];
                Memory[224]   <=  Memory[224];
                Memory[225]   <=  Memory[225];
                Memory[226]   <=  Memory[226];
                Memory[227]   <=  Memory[227];
                Memory[228]   <=  Memory[228];
                Memory[229]   <=  Memory[229];
                Memory[230]   <=  Memory[230];
                Memory[231]   <=  Memory[231];
                Memory[232]   <=  Memory[232];
                Memory[233]   <=  Memory[233];
                Memory[234]   <=  Memory[234];
                Memory[235]   <=  Memory[235];
                Memory[236]   <=  Memory[236];
                Memory[237]   <=  Memory[237];
                Memory[238]   <=  Memory[238];
                Memory[239]   <=  Memory[239];
                Memory[240]   <=  Memory[240];
                Memory[241]   <=  Memory[241];
                Memory[242]   <=  Memory[242];
                Memory[243]   <=  Memory[243];
                Memory[244]   <=  Memory[244];
                Memory[245]   <=  Memory[245];
                Memory[246]   <=  Memory[246];
                Memory[247]   <=  Memory[247];
                Memory[248]   <=  Memory[248];
                Memory[249]   <=  Memory[249];
                Memory[250]   <=  Memory[250];
                Memory[251]   <=  Memory[251];
                Memory[252]   <=  Memory[252];
                Memory[253]   <=  Memory[253];
                Memory[254]   <=  Memory[254];
                Memory[255]   <=  Memory[255];
            end
        end
    end
endmodule

